class apb_config_db;

static mailbox gen2bfm=new();
static mailbox mon2scb=new();
static virtual apb_interface cfg_intf_h;
endclass
